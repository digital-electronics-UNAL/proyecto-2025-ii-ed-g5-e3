module LCD1602_controllerP #(parameter NUM_COMMANDS = 4, 
                                      NUM_DATA_ALL = 32,  
                                      NUM_DATA_PERLINE = 16,
                                      DATA_BITS = 8,
                                      COUNT_MAX = 800000)(
    input clk,            
    input reset,          
    input ready_i,
    output reg rs,        
    output reg rw,
    output enable,    
    output reg [DATA_BITS-1:0] data
);

localparam IDLE = 3'b000;
localparam CONFIG_CMD1 = 3'b001;
localparam WR_STATIC_TEXT_1L = 3'b010;
localparam CONFIG_CMD2 = 3'b011;
localparam WR_STATIC_TEXT_2L = 3'b100;
localparam WR_Din_TEXT = 3'b101;

localparam SetCursor=2'b00;
localparam WR_Din_DATA=2'b01;
localparam SetCursor2=2'b10;
localparam WR_Din_DATA2=2'b11;

reg [2:0] fsm_state;
reg [2:0] next_state;
reg clk_16ms;
reg [1:0] sel_dinamic;

localparam CLEAR_DISPLAY = 8'h01;
localparam SHIFT_CURSOR_RIGHT = 8'h06;
localparam DISPON_CURSOROFF = 8'h0C;
localparam LINES2_MATRIX5x8_MODE8bit = 8'h38;
localparam START_2LINE = 8'hC0;

reg [$clog2(COUNT_MAX)-1:0] clk_counter;
reg [$clog2(NUM_COMMANDS):0] command_counter;
reg [$clog2(NUM_DATA_PERLINE):0] data_counter;

reg [DATA_BITS-1:0] static_data_mem [0: NUM_DATA_ALL-1];
reg [DATA_BITS-1:0] config_mem [0:NUM_COMMANDS-1]; 

reg [4:0] dot_count = 0;
reg [7:0] dot_mem [0:15];
reg [$clog2(16):0] i;

initial begin
    fsm_state <= IDLE;
    command_counter <= 'b0;
    data_counter <= 'b0;
    rs <= 1'b0;
    rw <= 1'b0;
    data <= 8'b0;
    clk_16ms <= 1'b0;
    clk_counter <= 'b0;
    $readmemh("/home/camilo/github-classroom/digital-electronics-UNAL/lab07-lcd-en-modo-paralelo-2025-ii-ed-g5-e3/src/data.txt", static_data_mem);    
    config_mem[0] <= LINES2_MATRIX5x8_MODE8bit;
    config_mem[1] <= SHIFT_CURSOR_RIGHT;
    config_mem[2] <= DISPON_CURSOROFF;
    config_mem[3] <= CLEAR_DISPLAY;
end

always @(posedge clk) begin
    if (clk_counter == COUNT_MAX-1) begin
        clk_16ms <= ~clk_16ms;
        clk_counter <= 'b0;
    end else begin
        clk_counter <= clk_counter + 1;
    end
end

always @(posedge clk_16ms)begin
    if(reset == 0)begin
        fsm_state <= IDLE;
    end else begin
        fsm_state <= next_state;
    end
end

always @(*) begin
    case(fsm_state)
        IDLE: begin
            next_state <= (ready_i)? CONFIG_CMD1 : IDLE;
        end
        CONFIG_CMD1: begin 
            next_state <= (command_counter == NUM_COMMANDS)? WR_STATIC_TEXT_1L : CONFIG_CMD1;
        end
        WR_STATIC_TEXT_1L: begin
            next_state <= (data_counter == NUM_DATA_PERLINE)? CONFIG_CMD2 : WR_STATIC_TEXT_1L;
        end
        CONFIG_CMD2: begin 
            next_state <= WR_STATIC_TEXT_2L;
        end
        WR_STATIC_TEXT_2L: begin
            next_state <= (data_counter == NUM_DATA_PERLINE)? WR_Din_TEXT : WR_STATIC_TEXT_2L;
        end
        WR_Din_TEXT: begin
            next_state <= WR_Din_TEXT;
        end
        default: next_state = IDLE;
    endcase
end

always @(posedge clk_16ms) begin
    if (reset == 0) begin
        command_counter <= 'b0;
        data_counter <= 'b0;
        data <= 'b0;
        $readmemh("/home/camilo/github-classroom/digital-electronics-UNAL/lab07-lcd-en-modo-paralelo-2025-ii-ed-g5-e3/src/data.txt", static_data_mem);
    end else begin
        case (next_state)
            IDLE: begin
                command_counter <= 'b0;
                data_counter <= 'b0;
                rs <= 1'b0;
                data  <= 'b0;
            end
            CONFIG_CMD1: begin
                rs <= 1'b0; 
                data <= config_mem[command_counter];
                command_counter <= command_counter + 1;
            end
            WR_STATIC_TEXT_1L: begin
                rs <= 1'b1; 
                data <= static_data_mem[data_counter];
                data_counter <= data_counter + 1;
            end
            CONFIG_CMD2: begin
                rs <= 1'b0; 
                data <= START_2LINE;
                data_counter <= 'b0;
            end
            WR_STATIC_TEXT_2L: begin
                rs <= 1'b1; 
                data <= static_data_mem[NUM_DATA_PERLINE + data_counter];
                data_counter <= data_counter + 1;
                sel_dinamic <= SetCursor2;
            end
            WR_Din_TEXT: begin
                case (sel_dinamic)
                    SetCursor2: begin
                        rs <= 1'b0;
                        data <= 8'hC0;   // cursor solo en la segunda línea
                        sel_dinamic <= WR_Din_DATA2;
                        data_counter <= 0;
                    end
                    WR_Din_DATA2: begin
                        rs <= 1'b1;
                        data <= dot_mem[data_counter];
                        if (data_counter == 15) begin
                            if (dot_count == 16)
                                dot_count <= 0;
                            else
                                dot_count <= dot_count + 1;
                            for (i = 0; i < 16; i = i + 1) begin
                                if (i < dot_count)
                                    dot_mem[i] <= 8'h2E;
                                else
                                    dot_mem[i] <= 8'h20;
                            end
                            sel_dinamic <= SetCursor2;
                        end else begin
                            data_counter <= data_counter + 1;
                            sel_dinamic <= WR_Din_DATA2;
                        end
                    end
                endcase
            end
        endcase
    end
end

assign enable = clk_16ms;

endmodule